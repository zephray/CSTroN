`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:53:22 08/16/2018 
// Design Name: 
// Module Name:    gldp_lut 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gldp_lut(
    input rst,
    input flm,
    input [4:0] raw_in,
    input inv,
    output reg dither_out
    );
    
    reg [31-1:0] gldp_lut_sr_a [0:31];
    reg [31-1:0] gldp_lut_sr_b [0:31];
    
    initial
    begin

        gldp_lut_sr_a[0]  = 31'b0000000000000000000000000000000;
        gldp_lut_sr_b[0]  = 31'b0000000000000000000000000000000;

        gldp_lut_sr_a[1]  = 31'b1000000000000000000000000000000;
        gldp_lut_sr_b[1]  = 31'b0000000000000001000000000000000;

        gldp_lut_sr_a[2]  = 31'b1000000000000001000000000000000;
        gldp_lut_sr_b[2]  = 31'b0000000100000000000000010000000;

        gldp_lut_sr_a[3]  = 31'b1000000000100000000001000000000;
        gldp_lut_sr_b[3]  = 31'b0000010000000001000000000100000;

        gldp_lut_sr_a[4]  = 31'b1000000010000000100000001000000;
        gldp_lut_sr_b[4]  = 31'b0000010000001000000010000000100;

        gldp_lut_sr_a[5]  = 31'b1000001000001000001000001000000;
        gldp_lut_sr_b[5]  = 31'b0010000010000001000001000001000;

        gldp_lut_sr_a[6]  = 31'b1000010000100001000010000100000;
        gldp_lut_sr_b[6]  = 31'b0010000100000100001000010000100;

        gldp_lut_sr_a[7]  = 31'b1000100001000100001000100001000;
        gldp_lut_sr_b[7]  = 31'b0010001000010001000100001000100;

        gldp_lut_sr_a[8]  = 31'b1000100010001000100010001000100;
        gldp_lut_sr_b[8]  = 31'b0010001000100010010001000100010;

        gldp_lut_sr_a[9]  = 31'b1001000100100010010001001000100;
        gldp_lut_sr_b[9]  = 31'b0100010010001001001000100100010;

        gldp_lut_sr_a[10] = 31'b1001001001001001001001001001000;
        gldp_lut_sr_b[10] = 31'b0100100100100010010010010010010;

        gldp_lut_sr_a[11] = 31'b1001001001001001001001001001001;
        gldp_lut_sr_b[11] = 31'b0100100100100110010010010010010;

        gldp_lut_sr_a[12] = 31'b1010010100101001001001010010100;
        gldp_lut_sr_b[12] = 31'b0100101001010010100101001010010;

        gldp_lut_sr_a[13] = 31'b1010100101010010101001010100100;
        gldp_lut_sr_b[13] = 31'b0101010010101001001010100101010;

        gldp_lut_sr_a[14] = 31'b1010101010010101010010101010100;
        gldp_lut_sr_b[14] = 31'b0101010010101010010101010100101;

        gldp_lut_sr_a[15] = 31'b1010101010101010101010101010100;
        gldp_lut_sr_b[15] = 31'b0101010101010100101010101010101;

        gldp_lut_sr_a[16] = 31'b0101010101010101010101010101011;
        gldp_lut_sr_b[16] = 31'b1010101010101011010101010101010;

        gldp_lut_sr_a[17] = 31'b0101010101101010101101010101011;
        gldp_lut_sr_b[17] = 31'b1010101101010101101010101011010;

        gldp_lut_sr_a[18] = 31'b0101011010101101010110101011011;
        gldp_lut_sr_b[18] = 31'b1010101101010110110101011010101;

        gldp_lut_sr_a[19] = 31'b0101101011010110110110101101011;
        gldp_lut_sr_b[19] = 31'b1011010110101101011010110101101;

        gldp_lut_sr_a[20] = 31'b0110110110110110110110110110110;
        gldp_lut_sr_b[20] = 31'b1011011011011001101101101101101;

        gldp_lut_sr_a[21] = 31'b0110110110110110110110110110111;
        gldp_lut_sr_b[21] = 31'b1011011011011101101101101101101;

        gldp_lut_sr_a[22] = 31'b0110111011011101101110110111011;
        gldp_lut_sr_b[22] = 31'b1011101101110110110111011011101;

        gldp_lut_sr_a[23] = 31'b0111011101110111011101110111011;
        gldp_lut_sr_b[23] = 31'b1101110111011101101110111011101;

        gldp_lut_sr_a[24] = 31'b0111011110111011110111011110111;
        gldp_lut_sr_b[24] = 31'b1101110111101110111011110111011;

        gldp_lut_sr_a[25] = 31'b0111101111011110111101111011111;
        gldp_lut_sr_b[25] = 31'b1101111011111011110111101111011;

        gldp_lut_sr_a[26] = 31'b0111110111110111110111110111111;
        gldp_lut_sr_b[26] = 31'b1101111101111110111110111110111;

        gldp_lut_sr_a[27] = 31'b0111111101111111011111110111111;
        gldp_lut_sr_b[27] = 31'b1111101111110111111101111111011;

        gldp_lut_sr_a[28] = 31'b0111111111011111111110111111111;
        gldp_lut_sr_b[28] = 31'b1111101111111110111111111011111;

        gldp_lut_sr_a[29] = 31'b0111111111111110111111111111111;
        gldp_lut_sr_b[29] = 31'b1111111011111111111111101111111;

        gldp_lut_sr_a[30] = 31'b0111111111111111111111111111111;
        gldp_lut_sr_b[30] = 31'b1111111111111110111111111111111;

        gldp_lut_sr_a[31] = 31'b1111111111111111111111111111111;
        gldp_lut_sr_b[31] = 31'b1111111111111111111111111111111;

    end
    
    
    integer i;
    
    always @(posedge flm, posedge rst)
    begin
        if (rst) begin
            // should we reset at all? Reset all SR to default value?
        end
        else begin
            for (i = 0; i < 32; i = i + 1) begin
                gldp_lut_sr_a[i] <= {gldp_lut_sr_a[i][29:0], gldp_lut_sr_a[i][30]};
                gldp_lut_sr_b[i] <= {gldp_lut_sr_b[i][29:0], gldp_lut_sr_b[i][30]};
            end
        end
    end
    
    always @(raw_in, inv) begin
        if (inv)
            dither_out = gldp_lut_sr_b[raw_in][0];
        else
            dither_out = gldp_lut_sr_a[raw_in][0];
    end

endmodule
