`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:53:22 08/16/2018 
// Design Name: 
// Module Name:    gldp_lut 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gldp_lut(
    input rst,
    input flm,
    input [4:0] raw_in,
    input inv,
    output reg dither_out
    );
    
    reg [49-1:0] gldp_lut_sr_a [0:31];
    reg [49-1:0] gldp_lut_sr_b [0:31];
    
    reg [5:0] gldp_inverse_counter = 0;
    reg       gldp_inverse_internal = 0;
    wire      gldp_inverse = gldp_inverse_internal ^ inv;
    
    initial
    begin
        gldp_lut_sr_a[0]  = 49'b0000000000000000000000000000000000000000000000000;
        gldp_lut_sr_b[0]  = 49'b0000000000000000000000000000000000000000000000000;

        gldp_lut_sr_a[1]  = 49'b0000000000000001000000000000000010000000000000001;
        gldp_lut_sr_b[1]  = 49'b0000000010000000000000001000000000000000100000000;

        gldp_lut_sr_a[2]  = 49'b0000000100000001000000010000000100000001000000001;
        gldp_lut_sr_b[2]  = 49'b0010000000100000000100000001000000010000000100000;

        gldp_lut_sr_a[3]  = 49'b0000001000000100000010000001000000100000010000001;
        gldp_lut_sr_b[3]  = 49'b0001000000100000010000001000000100000010000001000;

        gldp_lut_sr_a[4]  = 49'b0000010000010000010000010000010000010000010000001;
        gldp_lut_sr_b[4]  = 49'b0010000010000010000001000001000001000001000001000;

        gldp_lut_sr_a[5]  = 49'b0000100001000010000100001000010000100001000010001;
        gldp_lut_sr_b[5]  = 49'b0010000100001000010001000010000100001000010000100;

        gldp_lut_sr_a[6]  = 49'b0001000100010001000100010001000100010001000100001;
        gldp_lut_sr_b[6]  = 49'b0100010001000100010000100010001000100010001000100;

        gldp_lut_sr_a[7]  = 49'b0001001000100100010010001001000100100010010001001;
        gldp_lut_sr_b[7]  = 49'b0100010010001001000100100010010001001000100100010;

        gldp_lut_sr_a[8]  = 49'b0010010010001001001001000100100100100010010010001;
        gldp_lut_sr_b[8]  = 49'b1000100100100100010010010001001001001000100100100;

        gldp_lut_sr_a[9]  = 49'b0010010010010010010010010010010010010010010010001;
        gldp_lut_sr_b[9]  = 49'b1001001001001001001000100100100100100100100100100;

        gldp_lut_sr_a[10] = 49'b0100100101001001010010010100100101001001010010010;
        gldp_lut_sr_b[10] = 49'b1010010010100100101001001001001001010010010100100;

        gldp_lut_sr_a[11] = 49'b0100101001010010100101010010100101001010010100101;
        gldp_lut_sr_b[11] = 49'b1001010010101001010010100101001010010101001010010;

        gldp_lut_sr_a[12] = 49'b0101010100101010100101010101001010101001010101001;
        gldp_lut_sr_b[12] = 49'b1010010101010010101010100101010100101010100101010;

        gldp_lut_sr_a[13] = 49'b0101010101010100101010101010100101010101010101001;
        gldp_lut_sr_b[13] = 49'b1010100101010101010100101010101010101001010101010;

        gldp_lut_sr_a[14] = 49'b0101010101010101010101010101010101010101010101010;
        gldp_lut_sr_b[14] = 49'b1010101010101010101010100101010101010101010101010;

        gldp_lut_sr_a[15] = 49'b0101010101010101101010101010101011010101010101011;
        gldp_lut_sr_b[15] = 49'b1010101011010101010101010110101010101010110101010;

        gldp_lut_sr_a[16] = 49'b0101010101101010101101010101011010101011010101011;
        gldp_lut_sr_b[16] = 49'b1010110101010110101010101101010101101010101101010;

        gldp_lut_sr_a[17] = 49'b0101011010110101101011010101101011010110101101011;
        gldp_lut_sr_b[17] = 49'b1011010110101101011010101101011010110101101011010;

        gldp_lut_sr_a[18] = 49'b0110110110101101101101011011011010110110110101101;
        gldp_lut_sr_b[18] = 49'b1101101101011011011010110110110101101101101011010;

        gldp_lut_sr_a[19] = 49'b0110110110110110110110110110110110110110110110111;
        gldp_lut_sr_b[19] = 49'b1011011011011011011011011101101101101101101101101;

        gldp_lut_sr_a[20] = 49'b0111011011011011101101101101110110110110111011011;
        gldp_lut_sr_b[20] = 49'b1101110110110110111011011011101101101101110110110;

        gldp_lut_sr_a[21] = 49'b0111101110110111011101101110111011011101110110111;
        gldp_lut_sr_b[21] = 49'b1111011101101110111011011101110110111011101101110;

        gldp_lut_sr_a[22] = 49'b0111011101110111011101110111011101110111011101111;
        gldp_lut_sr_b[22] = 49'b1011101110111011101111011101110111011101110111011;

        gldp_lut_sr_a[23] = 49'b0111011110111011110111011110111011110111011110111;
        gldp_lut_sr_b[23] = 49'b1101110111101110111101110111011110111011110111011;

        gldp_lut_sr_a[24] = 49'b0111101111011110111101111011110111101111011110111;
        gldp_lut_sr_b[24] = 49'b1101111011110111101111011101111011110111101111011;

        gldp_lut_sr_a[25] = 49'b0111110111110111110111110111110111110111110111111;
        gldp_lut_sr_b[25] = 49'b1101111101111101111101111110111110111110111110111;

        gldp_lut_sr_a[26] = 49'b0111111011111101111110111111011111101111110111111;
        gldp_lut_sr_b[26] = 49'b1110111111011111101111110111111011111101111110111;

        gldp_lut_sr_a[27] = 49'b0111111101111111011111110111111101111111011111111;
        gldp_lut_sr_b[27] = 49'b1101111111011111110111111110111111101111111011111;

        gldp_lut_sr_a[28] = 49'b0111111111011111111101111111110111111111011111111;
        gldp_lut_sr_b[28] = 49'b1111101111111110111111110111111111011111111101111;

        gldp_lut_sr_a[29] = 49'b0111111111110111111111110111111111110111111111111;
        gldp_lut_sr_b[29] = 49'b1111111011111111111101111111111101111111111101111;

        gldp_lut_sr_a[30] = 49'b0111111111111111011111111111111101111111111111111;
        gldp_lut_sr_b[30] = 49'b1111111011111111111111110111111111111111011111111;

        gldp_lut_sr_a[31] = 49'b1111111111111111111111111111111111111111111111111;
        gldp_lut_sr_b[31] = 49'b1111111111111111111111111111111111111111111111111;
    end
    
    
    integer i;
    
    always @(posedge flm, posedge rst)
    begin
        if (rst) begin
            // should we reset at all? Reset all SR to default value?
        end
        else begin
            for (i = 0; i < 32; i = i + 1) begin
                gldp_lut_sr_a[i] <= {gldp_lut_sr_a[i][47:0], gldp_lut_sr_a[i][48]};
                gldp_lut_sr_b[i] <= {gldp_lut_sr_b[i][47:0], gldp_lut_sr_b[i][48]};
            end
            if (gldp_inverse_counter < (6'd49 - 1))
                gldp_inverse_counter <= gldp_inverse_counter + 1'b1;
            else begin
                gldp_inverse_counter <= 0;
                gldp_inverse_internal <= ~gldp_inverse_internal;
            end
        end
    end
    
    always @(raw_in, gldp_inverse) begin
        if (gldp_inverse)
            dither_out = gldp_lut_sr_b[raw_in][0];
        else
            dither_out = gldp_lut_sr_a[raw_in][0];
    end

endmodule
